library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

package my_types is
    type segment is (a,b,c,d,e);
end my_types;

package body my_types is
end my_types;